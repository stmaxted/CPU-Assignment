library IEEE;
use IEEE.std_logic_1164;
use IEEE.numeric_std.all;

entity CPU is
port (
			--Port Mapping here
		);
end entity CPU;


---------------------Functions to implement----------------------------
--		Conditional Branch
-- 	Unconditional Branch
--		Function Call (Jump)
--		Reading Data from memory
--		Writing data to memory
--		Arithmatic or Logic operation
-------------------------------------------------------------------------



architecture compute of CPU is
	--Aliases go here
begin

process(	--Sensitivity list) is
	--Variables
	begin
		--Outputs <= (others => '-');
		
	
	
	end process;
end architecture;